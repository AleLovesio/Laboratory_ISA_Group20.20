LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;


ENTITY abs_val IS
	GENERIC (N : INTEGER := 32);
	PORT (
		INPUT : IN SIGNED (N-1 DOWNTO 0);
		OUTPUT : OUT SIGNED (N-1 DOWNTO 0)); 
END ENTITY abs_val;

ARCHITECTURE UltraBehavioral OF abs_val IS
BEGIN  
	OUTPUT <= abs(INPUT);
END UltraBehavioral;

ARCHITECTURE Behavioral OF abs_val IS
SIGNAL COMPL_INPUT, NEG_OUTPUT : SIGNED (N-1 DOWNTO 0);
BEGIN  
	COMPL_INPUT <= NOT INPUT;
	NEG_OUTPUT <= COMPL_INPUT + 1;
	OUTPUT <= INPUT WHEN INPUT(N-1) = '0' ELSE NEG_OUTPUT;
END Behavioral;

ARCHITECTURE Behavioral_codelike OF abs_val IS
SIGNAL COMPL_INPUT, MSB_CIN, SIGN_VECT : SIGNED (N-1 DOWNTO 0);
BEGIN  
	SIGN_VECT <= SHIFT_RIGHT(INPUT, 31);
	COMPL_INPUT <= INPUT XOR SIGN_VECT;
	MSB_CIN <= TO_SIGNED(1, 32) AND SIGN_VECT;
	OUTPUT <= COMPL_INPUT + MSB_CIN;
END Behavioral_codelike;
