LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux2to1 IS
	GENERIC (N : INTEGER := 1); -- MUX X PARALLELISM
	PORT 	(	
				SEL		: IN STD_LOGIC; -- SELECTOR
				X0, X1	:IN STD_LOGIC_VECTOR (N-1 DOWNTO 0); -- INPUTS
				Y		: OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0) -- OUTPUT
			);
END ENTITY mux2to1;

ARCHITECTURE Behavioral OF mux2to1 IS
BEGIN
	Y <= X0 WHEN SEL = '0' ELSE X1;
END ARCHITECTURE Behavioral;