LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY imm_gen IS
	PORT(
			INSTRUCTION : IN STD_LOGIC_VECTOR (31 DOWNTO 0); 
			IMMEDIATE : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
		); 
END ENTITY imm_gen;

ARCHITECTURE Behavioral OF imm_gen IS
	--TYPE OPCODE IS (add, addi, auipc, lui, beq, lw, srai, andi, op_xor, slt, jal, sw) 
	-- ADD - R TYPE
	CONSTANT OPCODE_ADD 	: STD_LOGIC_VECTOR(6 DOWNTO 0)	:= "0110011";
	CONSTANT FUNCT3_ADD 	: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "000";
	-- ADDI - I TYPE
	CONSTANT OPCODE_ADDI 	: STD_LOGIC_VECTOR(6 DOWNTO 0)	:= "0010011";
	CONSTANT FUNCT3_ADDI 	: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "000";
	-- AUIPC - U TYPE
	CONSTANT OPCODE_AUIPC 	: STD_LOGIC_VECTOR(6 DOWNTO 0)	:= "0010111";
	-- LUI - U TYPE
	CONSTANT OPCODE_LUI 	: STD_LOGIC_VECTOR(6 DOWNTO 0)	:= "0110111";
	-- BEQ - B TYPE
	CONSTANT OPCODE_BEQ 	: STD_LOGIC_VECTOR(6 DOWNTO 0)	:= "1100011";
	CONSTANT FUNCT3_BEQ 	: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "000";
	-- LW - I TYPE
	CONSTANT OPCODE_LW 		: STD_LOGIC_VECTOR(6 DOWNTO 0)	:= "0000011";
	CONSTANT FUNCT3_LW 		: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "010";
	-- SRAI - R TYPE
	CONSTANT OPCODE_SRAI 	: STD_LOGIC_VECTOR(6 DOWNTO 0)	:= "0010011";
	CONSTANT FUNCT3_SRAI 	: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "101";
	-- ANDI - I TYPE
	CONSTANT OPCODE_ANDI 	: STD_LOGIC_VECTOR(6 DOWNTO 0) 	:= "0010011";
	CONSTANT FUNCT3_ANDI 	: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "111";
	-- XOR - R TYPE
	CONSTANT OPCODE_XOR 	: STD_LOGIC_VECTOR(6 DOWNTO 0) 	:= "0110011";
	CONSTANT FUNCT3_XOR 	: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "100";
	-- SLT - R TYPE
	CONSTANT OPCODE_SLT 	: STD_LOGIC_VECTOR(6 DOWNTO 0) 	:= "0110011";
	CONSTANT FUNCT3_SLT 	: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "010";
	-- JAL - J TYPE
	CONSTANT OPCODE_JAL 	: STD_LOGIC_VECTOR(6 DOWNTO 0)	:= "1101111";
	-- SW - S TYPE
	CONSTANT OPCODE_SW 		: STD_LOGIC_VECTOR(6 DOWNTO 0) 	:= "0100011";
	CONSTANT FUNCT3_SW	 	: STD_LOGIC_VECTOR(2 DOWNTO 0)	:= "010";
	
	CONSTANT ZEROS_31_0		: STD_LOGIC_VECTOR(31 DOWNTO 0)	:= (OTHERS => '0');
	CONSTANT ZEROS_11_0		: STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
	CONSTANT ZEROS_0		: STD_LOGIC						:= '0';
	
	SIGNAL 	 OPCODE			: STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL   FUNCT3			: STD_LOGIC_VECTOR(14 DOWNTO 12);
	SIGNAL	 R_TYPE_IMMEDIATE, I_TYPE_IMMEDIATE, S_TYPE_IMMEDIATE, B_TYPE_IMMEDIATE, U_TYPE_IMMEDIATE, J_TYPE_IMMEDIATE : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL   I_TYPE_IMMEDIATE_SHORT, S_TYPE_IMMEDIATE_SHORT : STD_LOGIC_VECTOR (11 DOWNTO 0); 
	SIGNAL   B_TYPE_IMMEDIATE_SHORT : STD_LOGIC_VECTOR (12 DOWNTO 0); 
	SIGNAL   J_TYPE_IMMEDIATE_SHORT : STD_LOGIC_VECTOR (20 DOWNTO 0);
	SIGNAL	 IS_R, IS_I, IS_S, IS_B, IS_U, IS_J : STD_LOGIC;
	
BEGIN
	OPCODE <= INSTRUCTION(6 DOWNTO 0);
	FUNCT3 <= INSTRUCTION(14 DOWNTO 12);
	
	I_TYPE_IMMEDIATE_SHORT <= INSTRUCTION(31 DOWNTO 20); 
	S_TYPE_IMMEDIATE_SHORT <= INSTRUCTION(31 DOWNTO 25) & INSTRUCTION(11 DOWNTO 7); 
	B_TYPE_IMMEDIATE_SHORT <= INSTRUCTION(31) & INSTRUCTION(7) & INSTRUCTION(30 DOWNTO 25) & INSTRUCTION(11 DOWNTO 8) & ZEROS_0; 
	J_TYPE_IMMEDIATE_SHORT <= INSTRUCTION(31) & INSTRUCTION(19 DOWNTO 12) & INSTRUCTION(20) & INSTRUCTION(30 DOWNTO 21) & ZEROS_0;
	
	R_TYPE_IMMEDIATE <= ZEROS_31_0;
	I_TYPE_IMMEDIATE <= STD_LOGIC_VECTOR(RESIZE(SIGNED(I_TYPE_IMMEDIATE_SHORT), I_TYPE_IMMEDIATE'LENGTH));
	S_TYPE_IMMEDIATE <= STD_LOGIC_VECTOR(RESIZE(SIGNED(S_TYPE_IMMEDIATE_SHORT), S_TYPE_IMMEDIATE'LENGTH));
	B_TYPE_IMMEDIATE <= STD_LOGIC_VECTOR(RESIZE(SIGNED(B_TYPE_IMMEDIATE_SHORT), B_TYPE_IMMEDIATE'LENGTH));
	U_TYPE_IMMEDIATE <= INSTRUCTION(31 DOWNTO 12) & ZEROS_11_0; 
	J_TYPE_IMMEDIATE <= STD_LOGIC_VECTOR(RESIZE(SIGNED(J_TYPE_IMMEDIATE_SHORT), J_TYPE_IMMEDIATE'LENGTH));
	
	IS_R <= '1' WHEN ((OPCODE = OPCODE_ADD) AND (FUNCT3 = FUNCT3_ADD)) OR ((OPCODE = OPCODE_SRAI) AND (FUNCT3 = FUNCT3_SRAI)) OR ((OPCODE = OPCODE_XOR) AND (FUNCT3 = FUNCT3_XOR)) OR ((OPCODE = OPCODE_SLT) AND (FUNCT3 = FUNCT3_SLT)) ELSE '0';
	IS_I <= '1' WHEN ((OPCODE = OPCODE_ADDI) AND (FUNCT3 = FUNCT3_ADDI)) OR ((OPCODE = OPCODE_LW) AND (FUNCT3 = FUNCT3_LW)) OR ((OPCODE = OPCODE_ANDI) AND (FUNCT3 = FUNCT3_ANDI)) ELSE '0';
	IS_S <= '1' WHEN ((OPCODE = OPCODE_SW) AND (FUNCT3 = FUNCT3_SW)) ELSE '0';
	IS_B <= '1' WHEN ((OPCODE = OPCODE_BEQ) AND (FUNCT3 = FUNCT3_BEQ)) ELSE '0';
	IS_U <= '1' WHEN (OPCODE = OPCODE_AUIPC) OR (OPCODE = OPCODE_LUI) ELSE '0';
	IS_J <= '1' WHEN (OPCODE = OPCODE_JAL) ELSE '0';
	
	IMMEDIATE <= 	R_TYPE_IMMEDIATE WHEN IS_R = '1' ELSE
					I_TYPE_IMMEDIATE WHEN IS_I = '1' ELSE
					S_TYPE_IMMEDIATE WHEN IS_S = '1' ELSE
					B_TYPE_IMMEDIATE WHEN IS_B = '1' ELSE
					U_TYPE_IMMEDIATE WHEN IS_U = '1' ELSE
					J_TYPE_IMMEDIATE WHEN IS_J = '1' ELSE
					ZEROS_31_0;
									
END ARCHITECTURE Behavioral;